module lut_ln 
#(
    parameter                           data_size = 32
)
(
    input                               clock_i                                                                 ,
    input                               reset_n_i                                                               ,
    input           [data_size/4 - 1:0] lut_ln_data_i                                                           ,
    input                               lut_ln_data_valid_i                                                     ,

    output                              lut_ln_data_valid_o                                                     ,
    output          [data_size - 1:0]   lut_ln_data_o
);
    integer                             i                                                                       ;
    reg             [data_size/2 - 1:0] LUT_LN  [255:0]                                                         ;

    reg             [data_size - 1:0]   lut_ln_data_o_temp                                                      ;
    reg                                 lut_ln_data_valid_o_temp                                                ;
    
    assign lut_ln_data_o = {lut_ln_data_o_temp, 16'b0}                                                          ;
    assign lut_ln_data_valid_o = lut_ln_data_valid_o_temp                                                       ;

    always @(posedge clock_i) 
    begin
        if (~reset_n_i)
            begin
                lut_ln_data_valid_o_temp <= 0                                                                   ;
                lut_ln_data_o_temp <= 0                                                                         ;
            end
        else
                if (lut_ln_data_valid_i && ~lut_ln_data_valid_o_temp)
                    begin
                        lut_ln_data_o_temp <= LUT_LN[lut_ln_data_i]                                             ;
                        lut_ln_data_valid_o_temp <= 1                                                           ;
                    end
    end


    //LUT LN (1,man) with man is 8 bits
    always @(posedge clock_i) 
    begin
        if (~reset_n_i)
            for (i = 0 ; i < 256 ; i = i + 1)
                LUT_LN[i] <= 0                                                                                  ;
        else
            begin
                LUT_LN[0] <= 16'b0000000000000000                                                               ;
                LUT_LN[1] <= 16'b0000000011111111                                                               ;
                LUT_LN[2] <= 16'b0000000111111110                                                               ;
                LUT_LN[3] <= 16'b0000001011111011                                                               ;
                LUT_LN[4] <= 16'b0000001111111000                                                               ;
                LUT_LN[5] <= 16'b0000010011110011                                                               ;
                LUT_LN[6] <= 16'b0000010111101110                                                               ;
                LUT_LN[7] <= 16'b0000011011100111                                                               ;
                LUT_LN[8] <= 16'b0000011111100000                                                               ;
                LUT_LN[9] <= 16'b0000100011011000                                                               ;
                LUT_LN[10] <= 16'b0000100111001111                                                              ;
                LUT_LN[11] <= 16'b0000101011000101                                                              ;
                LUT_LN[12] <= 16'b0000101110111010                                                              ;
                LUT_LN[13] <= 16'b0000110010101110                                                              ;
                LUT_LN[14] <= 16'b0000110110100001                                                              ;
                LUT_LN[15] <= 16'b0000111010010011                                                              ;
                LUT_LN[16] <= 16'b0000111110000101                                                              ;
                LUT_LN[17] <= 16'b0001000001110101                                                              ;
                LUT_LN[18] <= 16'b0001000101100101                                                              ;
                LUT_LN[19] <= 16'b0001001001010011                                                              ;
                LUT_LN[20] <= 16'b0001001101000001                                                              ;
                LUT_LN[21] <= 16'b0001010000101110                                                              ;
                LUT_LN[22] <= 16'b0001010100011011                                                              ;
                LUT_LN[23] <= 16'b0001011000000110                                                              ;
                LUT_LN[24] <= 16'b0001011011110000                                                              ;
                LUT_LN[25] <= 16'b0001011111011010                                                              ;
                LUT_LN[26] <= 16'b0001100011000011                                                              ;
                LUT_LN[27] <= 16'b0001100110101011                                                              ;
                LUT_LN[28] <= 16'b0001101010010010                                                              ;
                LUT_LN[29] <= 16'b0001101101111000                                                              ;
                LUT_LN[30] <= 16'b0001110001011110                                                              ;
                LUT_LN[31] <= 16'b0001110101000011                                                              ;
                LUT_LN[32] <= 16'b0001111000100111                                                              ;
                LUT_LN[33] <= 16'b0001111100001010                                                              ;
                LUT_LN[34] <= 16'b0001111111101100                                                              ;
                LUT_LN[35] <= 16'b0010000011001110                                                              ;
                LUT_LN[36] <= 16'b0010000110101110                                                              ;
                LUT_LN[37] <= 16'b0010001010001111                                                              ;
                LUT_LN[38] <= 16'b0010001101101110                                                              ;
                LUT_LN[39] <= 16'b0010010001001100                                                              ;
                LUT_LN[40] <= 16'b0010010100101010                                                              ;
                LUT_LN[41] <= 16'b0010011000000111                                                              ;
                LUT_LN[42] <= 16'b0010011011100011                                                              ;
                LUT_LN[43] <= 16'b0010011110111111                                                              ;
                LUT_LN[44] <= 16'b0010100010011010                                                              ;
                LUT_LN[45] <= 16'b0010100101110100                                                              ;
                LUT_LN[46] <= 16'b0010101001001101                                                              ;
                LUT_LN[47] <= 16'b0010101100100110                                                              ;
                LUT_LN[48] <= 16'b0010101111111110                                                              ;
                LUT_LN[49] <= 16'b0010110011010101                                                              ;
                LUT_LN[50] <= 16'b0010110110101100                                                              ;
                LUT_LN[51] <= 16'b0010111010000001                                                              ;
                LUT_LN[52] <= 16'b0010111101010111                                                              ;
                LUT_LN[53] <= 16'b0011000000101011                                                              ;
                LUT_LN[54] <= 16'b0011000011111111                                                              ;
                LUT_LN[55] <= 16'b0011000111010010                                                              ;
                LUT_LN[56] <= 16'b0011001010100100                                                              ;
                LUT_LN[57] <= 16'b0011001101110110                                                              ;
                LUT_LN[58] <= 16'b0011010001000111                                                              ;
                LUT_LN[59] <= 16'b0011010100010111                                                              ;
                LUT_LN[60] <= 16'b0011010111100111                                                              ;
                LUT_LN[61] <= 16'b0011011010110110                                                              ;
                LUT_LN[62] <= 16'b0011011110000101                                                              ;
                LUT_LN[63] <= 16'b0011100001010010                                                              ;
                LUT_LN[64] <= 16'b0011100100011111                                                              ;
                LUT_LN[65] <= 16'b0011100111101100                                                              ;
                LUT_LN[66] <= 16'b0011101010111000                                                              ;
                LUT_LN[67] <= 16'b0011101110000011                                                              ;
                LUT_LN[68] <= 16'b0011110001001110                                                              ;
                LUT_LN[69] <= 16'b0011110100011000                                                              ;
                LUT_LN[70] <= 16'b0011110111100001                                                              ;
                LUT_LN[71] <= 16'b0011111010101010                                                              ;
                LUT_LN[72] <= 16'b0011111101110010                                                              ;
                LUT_LN[73] <= 16'b0100000000111001                                                              ;
                LUT_LN[74] <= 16'b0100000100000000                                                              ;
                LUT_LN[75] <= 16'b0100000111000110                                                              ;
                LUT_LN[76] <= 16'b0100001010001100                                                              ;
                LUT_LN[77] <= 16'b0100001101010001                                                              ;
                LUT_LN[78] <= 16'b0100010000010110                                                              ;
                LUT_LN[79] <= 16'b0100010011011010                                                              ;
                LUT_LN[80] <= 16'b0100010110011101                                                              ;
                LUT_LN[81] <= 16'b0100011001100000                                                              ;
                LUT_LN[82] <= 16'b0100011100100010                                                              ;
                LUT_LN[83] <= 16'b0100011111100011                                                              ;
                LUT_LN[84] <= 16'b0100100010100101                                                              ;
                LUT_LN[85] <= 16'b0100100101100101                                                              ;
                LUT_LN[86] <= 16'b0100101000100101                                                              ;
                LUT_LN[87] <= 16'b0100101011100100                                                              ;
                LUT_LN[88] <= 16'b0100101110100011                                                              ;
                LUT_LN[89] <= 16'b0100110001100001                                                              ;
                LUT_LN[90] <= 16'b0100110100011111                                                              ;
                LUT_LN[91] <= 16'b0100110111011100                                                              ;
                LUT_LN[92] <= 16'b0100111010011001                                                              ;
                LUT_LN[93] <= 16'b0100111101010101                                                              ;
                LUT_LN[94] <= 16'b0101000000010000                                                              ;
                LUT_LN[95] <= 16'b0101000011001011                                                              ;
                LUT_LN[96] <= 16'b0101000110000110                                                              ;
                LUT_LN[97] <= 16'b0101001001000000                                                              ;
                LUT_LN[98] <= 16'b0101001011111001                                                              ;
                LUT_LN[99] <= 16'b0101001110110010                                                              ;
                LUT_LN[100] <= 16'b0101010001101010                                                             ;
                LUT_LN[101] <= 16'b0101010100100010                                                             ;
                LUT_LN[102] <= 16'b0101010111011001                                                             ;
                LUT_LN[103] <= 16'b0101011010010000                                                             ;
                LUT_LN[104] <= 16'b0101011101000110                                                             ;
                LUT_LN[105] <= 16'b0101011111111100                                                             ;
                LUT_LN[106] <= 16'b0101100010110010                                                             ;
                LUT_LN[107] <= 16'b0101100101100110                                                             ;
                LUT_LN[108] <= 16'b0101101000011011                                                             ;
                LUT_LN[109] <= 16'b0101101011001110                                                             ;
                LUT_LN[110] <= 16'b0101101110000010                                                             ;
                LUT_LN[111] <= 16'b0101110000110101                                                             ;
                LUT_LN[112] <= 16'b0101110011100111                                                             ;
                LUT_LN[113] <= 16'b0101110110011001                                                             ;
                LUT_LN[114] <= 16'b0101111001001010                                                             ;
                LUT_LN[115] <= 16'b0101111011111011                                                             ;
                LUT_LN[116] <= 16'b0101111110101011                                                             ;
                LUT_LN[117] <= 16'b0110000001011011                                                             ;
                LUT_LN[118] <= 16'b0110000100001011                                                             ;
                LUT_LN[119] <= 16'b0110000110111010                                                             ;
                LUT_LN[120] <= 16'b0110001001101000                                                             ;
                LUT_LN[121] <= 16'b0110001100010110                                                             ;
                LUT_LN[122] <= 16'b0110001111000100                                                             ;
                LUT_LN[123] <= 16'b0110010001110001                                                             ;
                LUT_LN[124] <= 16'b0110010100011110                                                             ;
                LUT_LN[125] <= 16'b0110010111001010                                                             ;
                LUT_LN[126] <= 16'b0110011001110110                                                             ;
                LUT_LN[127] <= 16'b0110011100100001                                                             ;
                LUT_LN[128] <= 16'b0110011111001100                                                             ;
                LUT_LN[129] <= 16'b0110100001110111                                                             ;
                LUT_LN[130] <= 16'b0110100100100001                                                             ;
                LUT_LN[131] <= 16'b0110100111001010                                                             ;
                LUT_LN[132] <= 16'b0110101001110011                                                             ;
                LUT_LN[133] <= 16'b0110101100011100                                                             ;
                LUT_LN[134] <= 16'b0110101111000100                                                             ;
                LUT_LN[135] <= 16'b0110110001101100                                                             ;
                LUT_LN[136] <= 16'b0110110100010011                                                             ;
                LUT_LN[137] <= 16'b0110110110111010                                                             ;
                LUT_LN[138] <= 16'b0110111001100001                                                             ;
                LUT_LN[139] <= 16'b0110111100000111                                                             ;
                LUT_LN[140] <= 16'b0110111110101101                                                             ;
                LUT_LN[141] <= 16'b0111000001010010                                                             ;
                LUT_LN[142] <= 16'b0111000011110111                                                             ;
                LUT_LN[143] <= 16'b0111000110011011                                                             ;
                LUT_LN[144] <= 16'b0111001000111111                                                             ;
                LUT_LN[145] <= 16'b0111001011100011                                                             ;
                LUT_LN[146] <= 16'b0111001110000110                                                             ;
                LUT_LN[147] <= 16'b0111010000101001                                                             ;
                LUT_LN[148] <= 16'b0111010011001011                                                             ;
                LUT_LN[149] <= 16'b0111010101101101                                                             ;
                LUT_LN[150] <= 16'b0111011000001111                                                             ;
                LUT_LN[151] <= 16'b0111011010110000                                                             ;
                LUT_LN[152] <= 16'b0111011101010001                                                             ;
                LUT_LN[153] <= 16'b0111011111110010                                                             ;
                LUT_LN[154] <= 16'b0111100010010010                                                             ;
                LUT_LN[155] <= 16'b0111100100110001                                                             ;
                LUT_LN[156] <= 16'b0111100111010001                                                             ;
                LUT_LN[157] <= 16'b0111101001101111                                                             ;
                LUT_LN[158] <= 16'b0111101100001110                                                             ;
                LUT_LN[159] <= 16'b0111101110101100                                                             ;
                LUT_LN[160] <= 16'b0111110001001010                                                             ;
                LUT_LN[161] <= 16'b0111110011100111                                                             ;
                LUT_LN[162] <= 16'b0111110110000100                                                             ;
                LUT_LN[163] <= 16'b0111111000100001                                                             ;
                LUT_LN[164] <= 16'b0111111010111101                                                             ;
                LUT_LN[165] <= 16'b0111111101011001                                                             ;
                LUT_LN[166] <= 16'b0111111111110100                                                             ;
                LUT_LN[167] <= 16'b1000000010001111                                                             ;
                LUT_LN[168] <= 16'b1000000100101010                                                             ;
                LUT_LN[169] <= 16'b1000000111000100                                                             ;
                LUT_LN[170] <= 16'b1000001001011110                                                             ;
                LUT_LN[171] <= 16'b1000001011111000                                                             ;
                LUT_LN[172] <= 16'b1000001110010001                                                             ;
                LUT_LN[173] <= 16'b1000010000101010                                                             ;
                LUT_LN[174] <= 16'b1000010011000011                                                             ;
                LUT_LN[175] <= 16'b1000010101011011                                                             ;
                LUT_LN[176] <= 16'b1000010111110011                                                             ;
                LUT_LN[177] <= 16'b1000011010001011                                                             ;
                LUT_LN[178] <= 16'b1000011100100010                                                             ;
                LUT_LN[179] <= 16'b1000011110111001                                                             ;
                LUT_LN[180] <= 16'b1000100001001111                                                             ;
                LUT_LN[181] <= 16'b1000100011100101                                                             ;
                LUT_LN[182] <= 16'b1000100101111011                                                             ;
                LUT_LN[183] <= 16'b1000101000010001                                                             ;
                LUT_LN[184] <= 16'b1000101010100110                                                             ;
                LUT_LN[185] <= 16'b1000101100111010                                                             ;
                LUT_LN[186] <= 16'b1000101111001111                                                             ;
                LUT_LN[187] <= 16'b1000110001100011                                                             ;
                LUT_LN[188] <= 16'b1000110011110111                                                             ;
                LUT_LN[189] <= 16'b1000110110001010                                                             ;
                LUT_LN[190] <= 16'b1000111000011101                                                             ;
                LUT_LN[191] <= 16'b1000111010110000                                                             ;
                LUT_LN[192] <= 16'b1000111101000010                                                             ;
                LUT_LN[193] <= 16'b1000111111010101                                                             ;
                LUT_LN[194] <= 16'b1001000001100110                                                             ;
                LUT_LN[195] <= 16'b1001000011111000                                                             ;
                LUT_LN[196] <= 16'b1001000110001001                                                             ;
                LUT_LN[197] <= 16'b1001001000011010                                                             ;
                LUT_LN[198] <= 16'b1001001010101010                                                             ;
                LUT_LN[199] <= 16'b1001001100111011                                                             ;
                LUT_LN[200] <= 16'b1001001111001010                                                             ;
                LUT_LN[201] <= 16'b1001010001011010                                                             ;
                LUT_LN[202] <= 16'b1001010011101001                                                             ;
                LUT_LN[203] <= 16'b1001010101111000                                                             ;
                LUT_LN[204] <= 16'b1001011000000111                                                             ;
                LUT_LN[205] <= 16'b1001011010010101                                                             ;
                LUT_LN[206] <= 16'b1001011100100011                                                             ;
                LUT_LN[207] <= 16'b1001011110110001                                                             ;
                LUT_LN[208] <= 16'b1001100000111110                                                             ;
                LUT_LN[209] <= 16'b1001100011001011                                                             ;
                LUT_LN[210] <= 16'b1001100101011000                                                             ;
                LUT_LN[211] <= 16'b1001100111100101                                                             ;
                LUT_LN[212] <= 16'b1001101001110001                                                             ;
                LUT_LN[213] <= 16'b1001101011111101                                                             ;
                LUT_LN[214] <= 16'b1001101110001000                                                             ;
                LUT_LN[215] <= 16'b1001110000010100                                                             ;
                LUT_LN[216] <= 16'b1001110010011111                                                             ;
                LUT_LN[217] <= 16'b1001110100101001                                                             ;
                LUT_LN[218] <= 16'b1001110110110100                                                             ;
                LUT_LN[219] <= 16'b1001111000111110                                                             ;
                LUT_LN[220] <= 16'b1001111011001000                                                             ;
                LUT_LN[221] <= 16'b1001111101010001                                                             ;
                LUT_LN[222] <= 16'b1001111111011010                                                             ;
                LUT_LN[223] <= 16'b1010000001100011                                                             ;
                LUT_LN[224] <= 16'b1010000011101100                                                             ;
                LUT_LN[225] <= 16'b1010000101110100                                                             ;
                LUT_LN[226] <= 16'b1010000111111100                                                             ;
                LUT_LN[227] <= 16'b1010001010000100                                                             ;
                LUT_LN[228] <= 16'b1010001100001100                                                             ;
                LUT_LN[229] <= 16'b1010001110010011                                                             ;
                LUT_LN[230] <= 16'b1010010000011010                                                             ;
                LUT_LN[231] <= 16'b1010010010100001                                                             ;
                LUT_LN[232] <= 16'b1010010100100111                                                             ;
                LUT_LN[233] <= 16'b1010010110101101                                                             ;
                LUT_LN[234] <= 16'b1010011000110011                                                             ;
                LUT_LN[235] <= 16'b1010011010111001                                                             ;
                LUT_LN[236] <= 16'b1010011100111110                                                             ;
                LUT_LN[237] <= 16'b1010011111000011                                                             ;
                LUT_LN[238] <= 16'b1010100001001000                                                             ;
                LUT_LN[239] <= 16'b1010100011001101                                                             ;
                LUT_LN[240] <= 16'b1010100101010001                                                             ;
                LUT_LN[241] <= 16'b1010100111010101                                                             ;
                LUT_LN[242] <= 16'b1010101001011001                                                             ;
                LUT_LN[243] <= 16'b1010101011011100                                                             ;
                LUT_LN[244] <= 16'b1010101101011111                                                             ;
                LUT_LN[245] <= 16'b1010101111100010                                                             ;
                LUT_LN[246] <= 16'b1010110001100101                                                             ;
                LUT_LN[247] <= 16'b1010110011100111                                                             ;
                LUT_LN[248] <= 16'b1010110101101010                                                             ;
                LUT_LN[249] <= 16'b1010110111101011                                                             ;
                LUT_LN[250] <= 16'b1010111001101101                                                             ;
                LUT_LN[251] <= 16'b1010111011101110                                                             ;
                LUT_LN[252] <= 16'b1010111101110000                                                             ;
                LUT_LN[253] <= 16'b1010111111110000                                                             ;
                LUT_LN[254] <= 16'b1011000001110001                                                             ;
                LUT_LN[255] <= 16'b1011000011110001                                                             ;
            end
    end
endmodule