/*
=====================================================================================
=                                                                                   =
=   Author: Hoang Van Quyen - UET - VNU                                             =
=                                                                                   =
=====================================================================================
*/
module lut_ln 
#(
    parameter                           data_size = 32
)
(
    input                               clock_i                                                                 ,
    input                               reset_n_i                                                               ,
    input           [data_size/4 - 1:0] lut_ln_data_i                                                           ,
    input                               lut_ln_data_valid_i                                                     ,

    output                              lut_ln_data_valid_o                                                     ,
    output          [data_size - 1:0]   lut_ln_data_o
);
    integer                             i                                                                       ;
    reg             [data_size - 1:0]   LUT_LN  [255:0]                                                         ;

    reg             [data_size - 1:0]   lut_ln_data_o_temp                                                      ;
    reg                                 lut_ln_data_valid_o_temp                                                ;
    
    assign lut_ln_data_o = lut_ln_data_o_temp                                                                   ;
    assign lut_ln_data_valid_o = lut_ln_data_valid_o_temp                                                       ;

    always @(posedge clock_i) 
    begin
        if (~reset_n_i)
            begin
                lut_ln_data_valid_o_temp <= 0                                                                   ;
                lut_ln_data_o_temp <= 0                                                                         ;
            end
        else
                if (lut_ln_data_valid_i && ~lut_ln_data_valid_o_temp)
                    begin
                        lut_ln_data_o_temp <= LUT_LN[lut_ln_data_i]                                             ;
                        lut_ln_data_valid_o_temp <= 1                                                           ;
                    end
    end


    //LUT LN (1,man) with man is 8 bits
    always @(posedge clock_i) 
    begin
        if (~reset_n_i)
            for (i = 0 ; i < 256 ; i = i + 1)
                LUT_LN[i] <= 0                                                                                  ;
        else
            begin
                LUT_LN[0]   <= 32'b00000000000000000000000000000000                                             ;
                LUT_LN[1]   <= 32'b00000000111111111000000001010101                                             ;
                LUT_LN[2]   <= 32'b00000001111111100000001010100110                                             ;
                LUT_LN[3]   <= 32'b00000010111110111000100011101100                                             ;
                LUT_LN[4]   <= 32'b00000011111110000001010100011000                                             ;
                LUT_LN[5]   <= 32'b00000100111100111010100100010000                                             ;
                LUT_LN[6]   <= 32'b00000101111011100100011011000000                                             ;
                LUT_LN[7]   <= 32'b00000110111001111111000000001000                                             ;
                LUT_LN[8]   <= 32'b00000111111000001010011011000000                                             ;
                LUT_LN[9]   <= 32'b00001000110110000110110011000000                                             ;
                LUT_LN[10]  <= 32'b00001001110011110100001111100000                                             ;
                LUT_LN[11]  <= 32'b00001010110001010010110111010000                                             ;
                LUT_LN[12]  <= 32'b00001011101110100010110010000000                                             ;
                LUT_LN[13]  <= 32'b00001100101011100100000110000000                                             ;
                LUT_LN[14]  <= 32'b00001101101000010110111011000000                                             ;
                LUT_LN[15]  <= 32'b00001110100100111011010111000000                                             ;
                LUT_LN[16]  <= 32'b00001111100001010001100001100000                                             ;
                LUT_LN[17]  <= 32'b00010000011101011001100001000000                                             ;
                LUT_LN[18]  <= 32'b00010001011001010011011011100000                                             ;
                LUT_LN[19]  <= 32'b00010010010100111111011000100000                                             ;
                LUT_LN[20]  <= 32'b00010011010000011101011110100000                                             ;
                LUT_LN[21]  <= 32'b00010100001011101101110011000000                                             ;
                LUT_LN[22]  <= 32'b00010101000110110000011101000000                                             ;
                LUT_LN[23]  <= 32'b00010110000001100101100010100000                                             ;
                LUT_LN[24]  <= 32'b00010110111100001101001010000000                                             ;
                LUT_LN[25]  <= 32'b00010111110110100111011001100000                                             ;
                LUT_LN[26]  <= 32'b00011000110000110100010111100000                                             ;
                LUT_LN[27]  <= 32'b00011001101010110100001001000000                                             ;
                LUT_LN[28]  <= 32'b00011010100100100110110101000000                                             ;
                LUT_LN[29]  <= 32'b00011011011110001100100000100000                                             ;
                LUT_LN[30]  <= 32'b00011100010111100101010010000000                                             ;
                LUT_LN[31]  <= 32'b00011101010000110001001111100000                                             ;
                LUT_LN[32]  <= 32'b00011110001001110000011101100000                                             ;
                LUT_LN[33]  <= 32'b00011111000010100011000011000000                                             ;
                LUT_LN[34]  <= 32'b00011111111011001001000101000000                                             ;
                LUT_LN[35]  <= 32'b00100000110011100010101001000000                                             ;
                LUT_LN[36]  <= 32'b00100001101011101111110100000000                                             ;
                LUT_LN[37]  <= 32'b00100010100011110000101100000000                                             ;
                LUT_LN[38]  <= 32'b00100011011011100101010111000000                                             ;
                LUT_LN[39]  <= 32'b00100100010011001101111001000000                                             ;
                LUT_LN[40]  <= 32'b00100101001010101010011000000000                                             ;
                LUT_LN[41]  <= 32'b00100110000001111010111001000000                                             ;
                LUT_LN[42]  <= 32'b00100110111000111111100001000000                                             ;
                LUT_LN[43]  <= 32'b00100111101111111000010110000000                                             ;
                LUT_LN[44]  <= 32'b00101000100110100101011011000000                                             ;
                LUT_LN[45]  <= 32'b00101001011101000110111000000000                                             ;
                LUT_LN[46]  <= 32'b00101010010011011100101111000000                                             ;
                LUT_LN[47]  <= 32'b00101011001001100111000111000000                                             ;
                LUT_LN[48]  <= 32'b00101011111111100110000100000000                                             ;
                LUT_LN[49]  <= 32'b00101100110101011001101010000000                                             ;
                LUT_LN[50]  <= 32'b00101101101011000001111111000000                                             ;
                LUT_LN[51]  <= 32'b00101110100000011111001000000000                                             ;
                LUT_LN[52]  <= 32'b00101111010101110001001000000000                                             ;
                LUT_LN[53]  <= 32'b00110000001010111000000101000000                                             ;
                LUT_LN[54]  <= 32'b00110000111111110100000011000000                                             ;
                LUT_LN[55]  <= 32'b00110001110100100101000111000000                                             ;
                LUT_LN[56]  <= 32'b00110010101001001011010101000000                                             ;
                LUT_LN[57]  <= 32'b00110011011101100110110001000000                                             ;
                LUT_LN[58]  <= 32'b00110100010001110111100001000000                                             ;
                LUT_LN[59]  <= 32'b00110101000101111101101000000000                                             ;
                LUT_LN[60]  <= 32'b00110101111001111001001010000000                                             ;
                LUT_LN[61]  <= 32'b00110110101101101010001101000000                                             ;
                LUT_LN[62]  <= 32'b00110111100001010000110100000000                                             ;
                LUT_LN[63]  <= 32'b00111000010100101101000011000000                                             ;
                LUT_LN[64]  <= 32'b00111001000111111110111110000000                                             ;
                LUT_LN[65]  <= 32'b00111001111011000110101010000000                                             ;
                LUT_LN[66]  <= 32'b00111010101110000100001011000000                                             ;
                LUT_LN[67]  <= 32'b00111011100000110111100101000000                                             ;
                LUT_LN[68]  <= 32'b00111100010011100000111011000000                                             ;
                LUT_LN[69]  <= 32'b00111101000110000000010011000000                                             ;
                LUT_LN[70]  <= 32'b00111101111000010101101110000000                                             ;
                LUT_LN[71]  <= 32'b00111110101010100001010011000000                                             ;
                LUT_LN[72]  <= 32'b00111111011100100011000011000000                                             ;
                LUT_LN[73]  <= 32'b01000000001110011011000100000000                                             ;
                LUT_LN[74]  <= 32'b01000001000000001001011010000000                                             ;
                LUT_LN[75]  <= 32'b01000001110001101110000110000000                                             ;
                LUT_LN[76]  <= 32'b01000010100011001001001110000000                                             ;
                LUT_LN[77]  <= 32'b01000011010100011010110110000000                                             ;
                LUT_LN[78]  <= 32'b01000100000101100011000000000000                                             ;
                LUT_LN[79]  <= 32'b01000100110110100001110000000000                                             ;
                LUT_LN[80]  <= 32'b01000101100111010111001010000000                                             ;
                LUT_LN[81]  <= 32'b01000110011000000011010010000000                                             ;
                LUT_LN[82]  <= 32'b01000111001000100110001100000000                                             ;
                LUT_LN[83]  <= 32'b01000111111000111111111010000000                                             ;
                LUT_LN[84]  <= 32'b01001000101001010000100000000000                                             ;
                LUT_LN[85]  <= 32'b01001001011001011000000010000000                                             ;
                LUT_LN[86]  <= 32'b01001010001001010110100010000000                                             ;
                LUT_LN[87]  <= 32'b01001010111001001100000100000000                                             ;
                LUT_LN[88]  <= 32'b01001011101000111000101100000000                                             ;
                LUT_LN[89]  <= 32'b01001100011000011100011100000000                                             ;
                LUT_LN[90]  <= 32'b01001101000111110111011010000000                                             ;
                LUT_LN[91]  <= 32'b01001101110111001001100110000000                                             ;
                LUT_LN[92]  <= 32'b01001110100110010011000110000000                                             ;
                LUT_LN[93]  <= 32'b01001111010101010011111010000000                                             ;
                LUT_LN[94]  <= 32'b01010000000100001100001000000000                                             ;
                LUT_LN[95]  <= 32'b01010000110010111011110010000000                                             ;
                LUT_LN[96]  <= 32'b01010001100001100010111100000000                                             ;
                LUT_LN[97]  <= 32'b01010010010000000001101000000000                                             ;
                LUT_LN[98]  <= 32'b01010010111110010111111010000000                                             ;
                LUT_LN[99]  <= 32'b01010011101100100101110100000000                                             ;
                LUT_LN[100] <= 32'b01010100011010101011011000000000                                             ;
                LUT_LN[101] <= 32'b01010101001000101000101100000000                                             ;
                LUT_LN[102] <= 32'b01010101110110011101110010000000                                             ;
                LUT_LN[103] <= 32'b01010110100100001010101100000000                                             ;
                LUT_LN[104] <= 32'b01010111010001101111011100000000                                             ;
                LUT_LN[105] <= 32'b01010111111111001100001000000000                                             ;
                LUT_LN[106] <= 32'b01011000101100100000110000000000                                             ;
                LUT_LN[107] <= 32'b01011001011001101101011000000000                                             ;
                LUT_LN[108] <= 32'b01011010000110110010000010000000                                             ;
                LUT_LN[109] <= 32'b01011010110011101110110010000000                                             ;
                LUT_LN[110] <= 32'b01011011100000100011101010000000                                             ;
                LUT_LN[111] <= 32'b01011100001101010000101110000000                                             ;
                LUT_LN[112] <= 32'b01011100111001110110000000000000                                             ;
                LUT_LN[113] <= 32'b01011101100110010011100010000000                                             ;
                LUT_LN[114] <= 32'b01011110010010101001010110000000                                             ;
                LUT_LN[115] <= 32'b01011110111110110111100000000000                                             ;
                LUT_LN[116] <= 32'b01011111101010111110000100000000                                             ;
                LUT_LN[117] <= 32'b01100000010110111101000010000000                                             ;
                LUT_LN[118] <= 32'b01100001000010110100011110000000                                             ;
                LUT_LN[119] <= 32'b01100001101110100100011010000000                                             ;
                LUT_LN[120] <= 32'b01100010011010001100111000000000                                             ;
                LUT_LN[121] <= 32'b01100011000101101101111100000000                                             ;
                LUT_LN[122] <= 32'b01100011110001000111101000000000                                             ;
                LUT_LN[123] <= 32'b01100100011100011001111110000000                                             ;
                LUT_LN[124] <= 32'b01100101000111100101000010000000                                             ;
                LUT_LN[125] <= 32'b01100101110010101000110100000000                                             ;
                LUT_LN[126] <= 32'b01100110011101100101011000000000                                             ;
                LUT_LN[127] <= 32'b01100111001000011010110000000000                                             ;
                LUT_LN[128] <= 32'b01100111110011001000111110000000                                             ;
                LUT_LN[129] <= 32'b01101000011101110000000110000000                                             ;
                LUT_LN[130] <= 32'b01101001001000010000001010000000                                             ;
                LUT_LN[131] <= 32'b01101001110010101001001010000000                                             ;
                LUT_LN[132] <= 32'b01101010011100111011001010000000                                             ;
                LUT_LN[133] <= 32'b01101011000111000110001100000000                                             ;
                LUT_LN[134] <= 32'b01101011110001001010010100000000                                             ;
                LUT_LN[135] <= 32'b01101100011011000111100000000000                                             ;
                LUT_LN[136] <= 32'b01101101000100111101111000000000                                             ;
                LUT_LN[137] <= 32'b01101101101110101101011010000000                                             ;
                LUT_LN[138] <= 32'b01101110011000010110001010000000                                             ;
                LUT_LN[139] <= 32'b01101111000001111000001000000000                                             ;
                LUT_LN[140] <= 32'b01101111101011010011011010000000                                             ;
                LUT_LN[141] <= 32'b01110000010100101000000000000000                                             ;
                LUT_LN[142] <= 32'b01110000111101110101111010000000                                             ;
                LUT_LN[143] <= 32'b01110001100110111101001110000000                                             ;
                LUT_LN[144] <= 32'b01110010001111111101111100000000                                             ;
                LUT_LN[145] <= 32'b01110010111000111000001000000000                                             ;
                LUT_LN[146] <= 32'b01110011100001101011110000000000                                             ;
                LUT_LN[147] <= 32'b01110100001010011000111010000000                                             ;
                LUT_LN[148] <= 32'b01110100110010111111101000000000                                             ;
                LUT_LN[149] <= 32'b01110101011011011111111010000000                                             ;
                LUT_LN[150] <= 32'b01110110000011111001110010000000                                             ;
                LUT_LN[151] <= 32'b01110110101100001101010100000000                                             ;
                LUT_LN[152] <= 32'b01110111010100011010100000000000                                             ;
                LUT_LN[153] <= 32'b01110111111100100001011010000000                                             ;
                LUT_LN[154] <= 32'b01111000100100100010000010000000                                             ;
                LUT_LN[155] <= 32'b01111001001100011100011010000000                                             ;
                LUT_LN[156] <= 32'b01111001110100010000100110000000                                             ;
                LUT_LN[157] <= 32'b01111010011011111110100110000000                                             ;
                LUT_LN[158] <= 32'b01111011000011100110011110000000                                             ;
                LUT_LN[159] <= 32'b01111011101011001000001100000000                                             ;
                LUT_LN[160] <= 32'b01111100010010100011110110000000                                             ;
                LUT_LN[161] <= 32'b01111100111001111001011100000000                                             ;
                LUT_LN[162] <= 32'b01111101100001001001000000000000                                             ;
                LUT_LN[163] <= 32'b01111110001000010010100100000000                                             ;
                LUT_LN[164] <= 32'b01111110101111010110001000000000                                             ;
                LUT_LN[165] <= 32'b01111111010110010011110010000000                                             ;
                LUT_LN[166] <= 32'b01111111111101001011100000000000                                             ;
                LUT_LN[167] <= 32'b10000000100011111101011000000000                                             ;
                LUT_LN[168] <= 32'b10000001001010101001010100000000                                             ;
                LUT_LN[169] <= 32'b10000001110001001111011100000000                                             ;
                LUT_LN[170] <= 32'b10000010010111101111110100000000                                             ;
                LUT_LN[171] <= 32'b10000010111110001010011000000000                                             ;
                LUT_LN[172] <= 32'b10000011100100011111001100000000                                             ;
                LUT_LN[173] <= 32'b10000100001010101110010000000000                                             ;
                LUT_LN[174] <= 32'b10000100110000110111101000000000                                             ;
                LUT_LN[175] <= 32'b10000101010110111011011000000000                                             ;
                LUT_LN[176] <= 32'b10000101111100111001011100000000                                             ;
                LUT_LN[177] <= 32'b10000110100010110001111000000000                                             ;
                LUT_LN[178] <= 32'b10000111001000100100110000000000                                             ;
                LUT_LN[179] <= 32'b10000111101110010010000100000000                                             ;
                LUT_LN[180] <= 32'b10001000010011111001110100000000                                             ;
                LUT_LN[181] <= 32'b10001000111001011100000100000000                                             ;
                LUT_LN[182] <= 32'b10001001011110111000110100000000                                             ;
                LUT_LN[183] <= 32'b10001010000100010000000100000000                                             ;
                LUT_LN[184] <= 32'b10001010101001100001111100000000                                             ;
                LUT_LN[185] <= 32'b10001011001110101110010100000000                                             ;
                LUT_LN[186] <= 32'b10001011110011110101011000000000                                             ;
                LUT_LN[187] <= 32'b10001100011000110111000000000000                                             ;
                LUT_LN[188] <= 32'b10001100111101110011011000000000                                             ;
                LUT_LN[189] <= 32'b10001101100010101010011000000000                                             ;
                LUT_LN[190] <= 32'b10001110000111011100000100000000                                             ;
                LUT_LN[191] <= 32'b10001110101100001000100000000000                                             ;
                LUT_LN[192] <= 32'b10001111010000101111101100000000                                             ;
                LUT_LN[193] <= 32'b10001111110101010001101000000000                                             ;
                LUT_LN[194] <= 32'b10010000011001101110011100000000                                             ;
                LUT_LN[195] <= 32'b10010000111110000110000000000000                                             ;
                LUT_LN[196] <= 32'b10010001100010011000011100000000                                             ;
                LUT_LN[197] <= 32'b10010010000110100101101100000000                                             ;
                LUT_LN[198] <= 32'b10010010101010101101111000000000                                             ;
                LUT_LN[199] <= 32'b10010011001110110001000000000000                                             ;
                LUT_LN[200] <= 32'b10010011110010101111000100000000                                             ;
                LUT_LN[201] <= 32'b10010100010110101000000000000000                                             ;
                LUT_LN[202] <= 32'b10010100111010011100000000000000                                             ;
                LUT_LN[203] <= 32'b10010101011110001011000000000000                                             ;
                LUT_LN[204] <= 32'b10010110000001110100111100000000                                             ;
                LUT_LN[205] <= 32'b10010110100101011010000000000000                                             ;
                LUT_LN[206] <= 32'b10010111001000111010001000000000                                             ;
                LUT_LN[207] <= 32'b10010111101100010101010100000000                                             ;
                LUT_LN[208] <= 32'b10011000001111101011101000000000                                             ;
                LUT_LN[209] <= 32'b10011000110010111101000000000000                                             ;
                LUT_LN[210] <= 32'b10011001010110001001101000000000                                             ;
                LUT_LN[211] <= 32'b10011001111001010001011000000000                                             ;
                LUT_LN[212] <= 32'b10011010011100010100010100000000                                             ;
                LUT_LN[213] <= 32'b10011010111111010010011100000000                                             ;
                LUT_LN[214] <= 32'b10011011100010001011111000000000                                             ;
                LUT_LN[215] <= 32'b10011100000101000000100000000000                                             ;
                LUT_LN[216] <= 32'b10011100100111110000011100000000                                             ;
                LUT_LN[217] <= 32'b10011101001010011011101000000000                                             ;
                LUT_LN[218] <= 32'b10011101101101000010001000000000                                             ;
                LUT_LN[219] <= 32'b10011110001111100100000000000000                                             ;
                LUT_LN[220] <= 32'b10011110110010000001001100000000                                             ;
                LUT_LN[221] <= 32'b10011111010100011001110100000000                                             ;
                LUT_LN[222] <= 32'b10011111110110101101110000000000                                             ;
                LUT_LN[223] <= 32'b10100000011000111101001000000000                                             ;
                LUT_LN[224] <= 32'b10100000111011000111111100000000                                             ;
                LUT_LN[225] <= 32'b10100001011101001110001100000000                                             ;
                LUT_LN[226] <= 32'b10100001111111001111111100000000                                             ;
                LUT_LN[227] <= 32'b10100010100001001101001100000000                                             ;
                LUT_LN[228] <= 32'b10100011000011000101111000000000                                             ;
                LUT_LN[229] <= 32'b10100011100100111010001000000000                                             ;
                LUT_LN[230] <= 32'b10100100000110101001111100000000                                             ;
                LUT_LN[231] <= 32'b10100100101000010101010000000000                                             ;
                LUT_LN[232] <= 32'b10100101001001111100001100000000                                             ;
                LUT_LN[233] <= 32'b10100101101011011110101100000000                                             ;
                LUT_LN[234] <= 32'b10100110001100111100110100000000                                             ;
                LUT_LN[235] <= 32'b10100110101110010110101000000000                                             ;
                LUT_LN[236] <= 32'b10100111001111101100000100000000                                             ;
                LUT_LN[237] <= 32'b10100111110000111101001000000000                                             ;
                LUT_LN[238] <= 32'b10101000010010001001111000000000                                             ;
                LUT_LN[239] <= 32'b10101000110011010010011000000000                                             ;
                LUT_LN[240] <= 32'b10101001010100010110100100000000                                             ;
                LUT_LN[241] <= 32'b10101001110101010110100000000000                                             ;
                LUT_LN[242] <= 32'b10101010010110010010001100000000                                             ;
                LUT_LN[243] <= 32'b10101010110111001001101100000000                                             ;
                LUT_LN[244] <= 32'b10101011010111111100111100000000                                             ;
                LUT_LN[245] <= 32'b10101011111000101100000000000000                                             ;
                LUT_LN[246] <= 32'b10101100011001010110111000000000                                             ;
                LUT_LN[247] <= 32'b10101100111001111101100100000000                                             ;
                LUT_LN[248] <= 32'b10101101011010100000001000000000                                             ;
                LUT_LN[249] <= 32'b10101101111010111110101000000000                                             ;
                LUT_LN[250] <= 32'b10101110011011011000111100000000                                             ;
                LUT_LN[251] <= 32'b10101110111011101111001100000000                                             ;
                LUT_LN[252] <= 32'b10101111011100000001010100000000                                             ;
                LUT_LN[253] <= 32'b10101111111100001111011100000000                                             ;
                LUT_LN[254] <= 32'b10110000011100011001100000000000                                             ;
                LUT_LN[255] <= 32'b10110000111100011111100000000000                                             ;
            end
    end
endmodule